`resetall
`timescale 1 ns / 1 ps
`default_nettype none

module EmuTrigger(
    input wire trigger
);

endmodule

`resetall
