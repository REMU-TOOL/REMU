`timescale 1 ns / 1 ps
`default_nettype none

module EmuClock (
    output wire clock
);

endmodule

`default_nettype wire
