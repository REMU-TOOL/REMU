`timescale 1ns / 1ps

`include "axi.vh"

module EmuTracePortImp #(
    parameter   DATA_WIDTH  = 1
)(
    input  wire                     clk,
    input  wire [DATA_WIDTH-1:0]    data
);

endmodule
