`timescale 1 ns / 1 ps
`default_nettype none

(* keep, emulib_component = "trigger" *)
module EmuTrigger(
    input trigger
);

endmodule
