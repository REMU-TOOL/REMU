`timescale 1 ns / 1 ps

module chain(
    (* __emu_extern_intf = "test" *)
    input                   ren1,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           raddr1,
    (* __emu_extern_intf = "test" *)
    output  [31:0]          rdata1,
    (* __emu_extern_intf = "test" *)
    input                   wen1,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           waddr1,
    (* __emu_extern_intf = "test" *)
    input   [31:0]          wdata1,
    (* __emu_extern_intf = "test" *)
    input                   ren2,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           raddr2,
    (* __emu_extern_intf = "test" *)
    output  [63:0]          rdata2,
    (* __emu_extern_intf = "test" *)
    input                   wen2,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           waddr2,
    (* __emu_extern_intf = "test" *)
    input   [63:0]          wdata2,
    (* __emu_extern_intf = "test" *)
    input                   ren3,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           raddr3,
    (* __emu_extern_intf = "test" *)
    output  [127:0]          rdata3,
    (* __emu_extern_intf = "test" *)
    input                   wen3,
    (* __emu_extern_intf = "test" *)
    input   [2:0]           waddr3,
    (* __emu_extern_intf = "test" *)
    input   [127:0]          wdata3
);

    wire clk;
    EmuClock clock(.clock(clk));

    mem #(
        .WIDTH(32),
        .DEPTH(8),
        .OFFSET(0),
        .SYNCREAD(1)
    )
    u_mem1 (
        .clk(clk),
        .ren(ren1),
        .raddr(raddr1),
        .rdata(rdata1),
        .wen(wen1),
        .waddr(waddr1),
        .wdata(wdata1)
    );

    mem #(
        .WIDTH(64),
        .DEPTH(8),
        .OFFSET(0),
        .SYNCREAD(1)
    )
    u_mem2 (
        .clk(clk),
        .ren(ren2),
        .raddr(raddr2),
        .rdata(rdata2),
        .wen(wen2),
        .waddr(waddr2),
        .wdata(wdata2)
    );

    mem #(
        .WIDTH(128),
        .DEPTH(8),
        .OFFSET(0),
        .SYNCREAD(1)
    )
    u_mem3 (
        .clk(clk),
        .ren(ren3),
        .raddr(raddr3),
        .rdata(rdata3),
        .wen(wen3),
        .waddr(waddr3),
        .wdata(wdata3)
    );

endmodule
