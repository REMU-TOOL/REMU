`timescale 1ns / 1ps

module test(

    input                       clk,
    input                       resetn,

    output                      trig,

    output reg                  pause,
    input                       do_pause,
    input                       do_resume,

    input                       ff_scan,
    input                       ff_dir,
    input   [63:0]              ff_sdi,
    output  [63:0]              ff_sdo,
    input                       ram_scan,
    input                       ram_dir,
    input   [63:0]              ram_sdi,
    output  [63:0]              ram_sdo,

    input                       up_req,
    input                       down_req,
    output                      up,
    output                      down,

    // for testbench use
    output                      dut_clk,

    output reg  [63:0]          count,
    input                       count_write,
    input   [63:0]              count_wdata,

    input                       step_write,
    input   [63:0]              step_wdata,
    output                      step_trig

);

    //reg clk = 0, rst = 1;
    wire rst = !resetn;
    //reg pause = 0;
    //reg ff_scan = 0, ff_dir = 0;
    //reg [63:0] ff_sdi = 0;
    //wire [63:0] ff_sdo;
    //reg ram_scan = 0, ram_dir = 0;
    //reg [63:0] ram_sdi = 0;
    //wire [63:0] ram_sdo;

    wire dut_stall;

    wire dut_clk, dut_clk_en;
    ClockGate clk_gate(
        .CLK(clk),
        .EN(dut_clk_en),
        .GCLK(dut_clk)
    );

    wire emu_dut_ff_clk, emu_dut_ff_clk_en;
    ClockGate dut_ff_clk_gate(
        .CLK(clk),
        .EN(emu_dut_ff_clk_en),
        .GCLK(emu_dut_ff_clk)
    );

    wire emu_dut_ram_clk, emu_dut_ram_clk_en;
    ClockGate dut_ram_clk_gate(
        .CLK(clk),
        .EN(emu_dut_ram_clk_en),
        .GCLK(emu_dut_ram_clk)
    );

    wire              mem_axi_awvalid;
	wire              mem_axi_awready;
	wire       [31:0] mem_axi_awaddr;

	wire              mem_axi_wvalid;
	wire              mem_axi_wready;
	wire       [31:0] mem_axi_wdata;
	wire       [ 3:0] mem_axi_wstrb;

	wire              mem_axi_bvalid;
	wire              mem_axi_bready;

	wire              mem_axi_arvalid;
	wire              mem_axi_arready;
	wire       [31:0] mem_axi_araddr;

	wire              mem_axi_rvalid;
	wire              mem_axi_rready;
	wire       [31:0] mem_axi_rdata;

    wire putchar_valid, putchar_ready;
    wire [7:0] putchar_data;

    assign putchar_ready = 1'b1;

    always @(posedge clk)
        if (dut_clk_en && putchar_valid)
            $write("%c", putchar_data);

    EMU_DUT emu_dut(
        .emu_clk            (clk),
        .emu_rst            (rst),
        .emu_ff_se          (ff_scan),
        .emu_ff_di          (ff_dir ? ff_sdi : ff_sdo),
        .emu_ff_do          (ff_sdo),
        .emu_ram_se         (ram_scan),
        .emu_ram_sd         (ram_dir),
        .emu_ram_di         (ram_sdi),
        .emu_ram_do         (ram_sdo),
        .emu_dut_ff_clk     (emu_dut_ff_clk),
        .emu_dut_ram_clk    (emu_dut_ram_clk),
        .emu_dut_rst        (rst),
        .emu_dut_trig       (trig),
        .emu_stall          (pause || dut_stall),
        .emu_stall_gen      (dut_stall),
        .emu_up_req         (up_req),
        .emu_down_req       (down_req),
        .emu_up_stat        (up),
        .emu_down_stat      (down),
        .emu_auto_0_dram_awvalid        (mem_axi_awvalid),
        .emu_auto_0_dram_awready        (mem_axi_awready),
        .emu_auto_0_dram_awaddr         (mem_axi_awaddr),
        .emu_auto_0_dram_awid           (),
        .emu_auto_0_dram_awlen          (),
        .emu_auto_0_dram_awsize         (),
        .emu_auto_0_dram_awburst        (),
        .emu_auto_0_dram_awlock         (),
        .emu_auto_0_dram_awcache        (),
        .emu_auto_0_dram_awprot         (),
        .emu_auto_0_dram_awqos          (),
        .emu_auto_0_dram_awregion       (),
        .emu_auto_0_dram_wvalid         (mem_axi_wvalid),
        .emu_auto_0_dram_wready         (mem_axi_wready),
        .emu_auto_0_dram_wdata          (mem_axi_wdata),
        .emu_auto_0_dram_wstrb          (mem_axi_wstrb),
        .emu_auto_0_dram_wlast          (),
        .emu_auto_0_dram_bvalid         (mem_axi_bvalid),
        .emu_auto_0_dram_bready         (mem_axi_bready),
        .emu_auto_0_dram_bresp          (2'b00),
        .emu_auto_0_dram_bid            (1'd0),
        .emu_auto_0_dram_arvalid        (mem_axi_arvalid),
        .emu_auto_0_dram_arready        (mem_axi_arready),
        .emu_auto_0_dram_araddr         (mem_axi_araddr),
        .emu_auto_0_dram_arid           (),
        .emu_auto_0_dram_arlen          (),
        .emu_auto_0_dram_arsize         (),
        .emu_auto_0_dram_arburst        (),
        .emu_auto_0_dram_arlock         (),
        .emu_auto_0_dram_arcache        (),
        .emu_auto_0_dram_arprot         (),
        .emu_auto_0_dram_arqos          (),
        .emu_auto_0_dram_arregion       (),
        .emu_auto_0_dram_rvalid         (mem_axi_rvalid),
        .emu_auto_0_dram_rready         (mem_axi_rready),
        .emu_auto_0_dram_rdata          (mem_axi_rdata),
        .emu_auto_0_dram_rresp          (2'b00),
        .emu_auto_0_dram_rid            (1'd0),
        .emu_auto_0_dram_rlast          (1'b1),
        .emu_putchar_valid              (putchar_valid),
        .emu_putchar_ready              (putchar_ready),
        .emu_putchar_data               (putchar_data)
    );

    reg [7:0] mem [0:64*1024-1];

    reg [31:0] reg_write_addr;
    reg [31:0] reg_write_data;
    reg [3:0] reg_write_strb;
    reg reg_write_addr_valid, reg_write_data_valid, reg_write_resp_valid;
    wire reg_write_addr_data_ok = reg_write_addr_valid && reg_write_data_valid;

    always @(posedge clk) begin
        if (rst) begin
            reg_write_addr          <= 12'd0;
            reg_write_data          <= 32'd0;
            reg_write_strb          <= 4'd0;
            reg_write_addr_valid    <= 1'b0;
            reg_write_data_valid    <= 1'b0;
            reg_write_resp_valid    <= 1'b0;
        end
        else begin
            if (mem_axi_awvalid && mem_axi_awready) begin
                reg_write_addr          <= mem_axi_awaddr;
                reg_write_addr_valid    <= 1'b1;
            end
            if (mem_axi_wvalid && mem_axi_wready) begin
                reg_write_data          <= mem_axi_wdata;
                reg_write_strb          <= mem_axi_wstrb;
                reg_write_data_valid    <= 1'b1;
            end
            if (reg_write_addr_data_ok) begin
                reg_write_addr_valid    <= 1'b0;
                reg_write_data_valid    <= 1'b0;
                reg_write_resp_valid    <= 1'b1;
            end
            if (mem_axi_bvalid && mem_axi_bready) begin
                reg_write_resp_valid    <= 1'b0;
            end
        end
    end

    always @(posedge clk) begin
        if (reg_write_addr_data_ok) begin
            if (reg_write_strb[0]) mem[reg_write_addr + 0] <= reg_write_data[ 7: 0];
            if (reg_write_strb[1]) mem[reg_write_addr + 1] <= reg_write_data[15: 8];
            if (reg_write_strb[2]) mem[reg_write_addr + 2] <= reg_write_data[23:16];
            if (reg_write_strb[3]) mem[reg_write_addr + 3] <= reg_write_data[31:24];
        end
    end

    assign mem_axi_awready    = !reg_write_addr_valid && !reg_write_resp_valid;
    assign mem_axi_wready     = !reg_write_data_valid;
    assign mem_axi_bvalid     = reg_write_resp_valid;

    reg [31:0] reg_read_addr;
    reg [31:0] reg_read_data;
    reg reg_read_addr_valid, reg_read_data_valid;
    wire reg_do_read = reg_read_addr_valid && !reg_read_data_valid;

    always @(posedge clk) begin
        if (rst) begin
            reg_read_addr       <= 12'd0;
            reg_read_data       <= 32'd0;
            reg_read_addr_valid <= 1'b0;
            reg_read_data_valid <= 1'b0;
        end
        else begin
            if (mem_axi_arvalid && mem_axi_arready) begin
                reg_read_addr       <= mem_axi_araddr;
                reg_read_addr_valid <= 1'b1;
            end
            if (reg_do_read) begin
                reg_read_data[ 7: 0] <= mem[reg_read_addr + 0];
                reg_read_data[15: 8] <= mem[reg_read_addr + 1];
                reg_read_data[23:16] <= mem[reg_read_addr + 2];
                reg_read_data[31:24] <= mem[reg_read_addr + 3];
                reg_read_data_valid <= 1'b1;
            end
            if (mem_axi_rvalid && mem_axi_rready) begin
                reg_read_addr_valid <= 1'b0;
                reg_read_data_valid <= 1'b0;
            end
        end
    end

    assign mem_axi_arready    = !reg_read_addr_valid;
    assign mem_axi_rvalid     = reg_read_data_valid;
    assign mem_axi_rdata      = reg_read_data;

    assign dut_clk_en = !pause && !dut_stall;
    assign emu_dut_ff_clk_en = !pause && !dut_stall || ff_scan;
    assign emu_dut_ram_clk_en = !pause && !dut_stall || ram_scan;

    initial begin
        if ($test$plusargs("DUMP")) begin
            $dumpfile(`DUMPFILE);
            $dumpvars();
        end
    end

    initial $readmemh("../../../design/picorv32/baremetal.hex", mem);

    always @(posedge clk)
        if (!resetn)
            count <= 64'd0;
        else if (count_write)
            count <= count_wdata;
        else if (dut_clk_en)
            count <= count + 64'd1;

    reg [63:0] step, step_next;

    always @(posedge clk)
        if (!resetn)
            step <= 64'd0;
        else
            step <= step_next;

    always @*
        if (step_write)
            step_next = step_wdata;
        else if (step == 64'd0)
            step_next = 64'd0;
        else if (dut_clk_en)
            step_next = step - 64'd1;

    assign step_trig = step != 64'd0 && step_next == 64'd0;

    always @(posedge clk)
        if (!resetn)
            pause <= 1'b0;
        else if (trig || step_trig || do_pause)
            pause <= 1'b1;
        else if (do_resume)
            pause <= 1'b0;

endmodule
