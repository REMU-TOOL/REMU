`timescale 1 ns / 1 ps
`default_nettype none

(* keep, noblackbox *)
module EmuReset (
    (* __emu_user_rst *)
    output wire reset
);

endmodule

`default_nettype wire
