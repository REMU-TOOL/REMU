`timescale 1 ns / 1 ps
`default_nettype none

module EmuTrigger #(
    parameter DESC = "<empty>"
)(
    input wire trigger
);

endmodule

`default_nettype wire
