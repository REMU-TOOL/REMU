`timescale 1 ns / 1 ps

(* emulib_reset *)
module EmuReset #(
    parameter DURATION_CYCLES = 100
)
(
    input clock,
    output reset
);

endmodule
