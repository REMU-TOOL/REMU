`timescale 1ns / 1ps
`default_nettype none

(* keep, noblackbox *)
module EmuClock (
    (* __emu_user_clk *)
    output wire clock
);

endmodule

`default_nettype wire
