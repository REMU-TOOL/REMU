`timescale 1 ns / 1 ps

(* emulib_clock *)
module EmuClock #(
    parameter FREQUENCY_MHZ = 100
)
(
    output clock
);

endmodule
