`timescale 1 ns / 1 ps

(* emulib_reset *)
module EmuReset #(
    parameter DURATION_NS = 100
)
(
    output reset
);

endmodule
