`timescale 1 ns / 1 ps

(* emulib_trigger *)
module EmuTrigger(
    input trigger
);

endmodule
