`timescale 1 ns / 1 ps

(* keep *)
module EmuTrigger #(
    parameter DESC = "<empty>"
)(
    input wire trigger
);

endmodule
