`timescale 1 ns / 1 ps

(* keep *)
module EmuTriggerImp #(
    parameter DESC = "<empty>"
)(
    input wire trigger
);

endmodule
