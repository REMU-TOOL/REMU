`timescale 1ns / 1ps

(* keep, noblackbox *)
module EmuClock (
    (* __emu_user_clk *)
    output wire clock
);

endmodule
