`timescale 1 ns / 1 ps

(* keep, emulib_component = "trigger" *)
module EmuTrigger(
    input trigger
);

endmodule
