`timescale 1 ns / 1 ps

(* keep, noblackbox *)
module EmuReset (
    (* __emu_user_rst *)
    output wire reset
);

endmodule
