`timescale 1 ns / 1 ps

(* keep, noblackbox *)
module EmuTrigger #(
    parameter DESC = "<empty>"
)(
    (* __emu_user_trig, __emu_user_trig_desc = DESC *)
    input wire trigger
);

endmodule
