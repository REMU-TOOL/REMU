`timescale 1 ns / 1 ps

(* keep *)
module EmuReset (
    output wire reset
);

endmodule
