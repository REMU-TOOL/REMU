`timescale 1ns / 1ps

(* keep, emulib_component = "putchar" *)
module PutCharDevice (
    input           clk,
    input           valid,
    input   [7:0]   data
);

endmodule
