`timescale 1 ns / 1 ps

(* keep *)
module EmuClock (
    output wire clock
);

endmodule
