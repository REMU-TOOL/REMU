`timescale 1 ns / 1 ps
`default_nettype none

(* keep *)
module EmuReset (
    output wire reset
);

endmodule

`default_nettype wire
