`timescale 1 ns / 1 ps

(* emulib_component = "trigger" *)
module EmuTrigger(
    input trigger
);

endmodule
