`define EMU_STAT                12'h000
`define EMU_CTRL                12'h004
`define EMU_CYCLE_LO            12'h008
`define EMU_CYCLE_HI            12'h00c
`define EMU_STEP                12'H010
`define EMU_DMA_RD_ADDR_LO      12'h020
`define EMU_DMA_RD_ADDR_HI      12'h024
`define EMU_DMA_RD_LEN          12'h028
`define EMU_DMA_RD_CSR          12'h02c
`define EMU_DMA_WR_ADDR_LO      12'h030
`define EMU_DMA_WR_ADDR_HI      12'h034
`define EMU_DMA_WR_LEN          12'h038
`define EMU_DMA_WR_CSR          12'h03c
